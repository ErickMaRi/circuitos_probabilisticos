WEIN OSCILATOR
.SUBCKT OPA132_0    1 2 3 4 5
*
C1   11 12 3.240E-12
C2    6  7 8.000E-12
CSS  10 99 1.000E-30
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
FB    7 99 POLY(5) VB VC VE VLP VLN 0 248.0E6 -250E6 250E6 250E6 -250E6
GA    6  0 11 12 402.0E-6
GCM   0  6 10 99 4.020E-9
ISS   3 10 DC 160.0E-6
HLIM 90  0 VLIM 1E3
J1   11  2 10 JX
J2   12  1 10 JX
R2    6  9 100.0E3
RD1   4 11 2.490E3
RD2   4 12 2.490E3
RO1   8  5 20
RO2   7 99 20
RP    3  4 7.500E3
RSS  10 99 1.250E6
VB    9  0 DC 0
VC    3 53 DC 1.200
VE   54  4 DC .9
VLIM  7  8 DC 0
VLP  91  0 DC 40
VLN   0 92 DC 40
.MODEL DX D(IS=800.0E-18)
.MODEL JX PJF(IS=2.500E-15 BETA=1.010E-3 VTO=-1)
.ENDS

.TEMP 27
.TRAN 15U 30M UIC

.OPTIONS ABSTOL=1U ITL2=200 TRTOL=1
.PROBE V(7,0)

VNeg        0 5 15
VPos        4 0 15
XU1         2 3 4 5 1 OPA132_0
DZ2         6 7  D_BZV80_1 
DZ1         6 8  D_BZV80_1 
R2          8 1 6K ; *DIST: UNIFORM 0 *
R5          7 3 800 ; *DIST: UNIFORM 0 * 
R4          0 7 200 ; *DIST: UNIFORM 0 * 
R3          3 1 2.08K ; *DIST: UNIFORM 0 * 
C1          9 1 10N IC=0 ; *DIST: NORMAL 0.05 * 
C2        4 2 10N IC=0 ; *DIST: NORMAL 0.05 *
R1          0 2 15K ; *DIST: UNIFORM 0 *
R6        2 9 15K ; *DIST: UNIFORM 0 *

.MODEL D_BZV80_1 D( IS=12.4F N=1 BV=6.2 IBV=7.5M RS=2.03 
+      CJO=30P VJ=683M M=315M FC=500M TT=25.9N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

.END
