LINEAL (PSpice format)
.TEMP 27
.TRAN 20N 10U

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V(4,0)

VIN         3 0 DC 0 AC 1 0
+ PULSE ( 0 1 0  0  0  1e19 1e20 )
R2 1 0 982.1674139468827
L2 2 1 988.5822310855177u IC=0
R1 3 2 1.0240122108546599K
lin         4 3 1M IC=0 
C1 4 2 1.029459944017509u

.END
