LEAKY INTEGRATE AND FIRE
.SUBCKT STDOPAMP  INP INM VP VM OUT
+ PARAMS: GAIN=200K RIN=2MEG RINC=1E9 ROUT=75 SLEWRATE=500K FPOLE1=5 FPOLE2=1MEG 
+         VDROPOH=1.9 VDROPOL=1.9 VOFFS=1M IBIAS=80N IOFFS=20N 
.PARAM PI = 3.141592
.PARAM IS = 1.0E-12
.PARAM VT = 0.02585
.PARAM IMAX = 100.0E-2
.PARAM C1 = {IMAX/SLEWRATE}
.PARAM R1 = {1/(2*PI*C1*FPOLE1)}
.PARAM GM1 = {GAIN/R1}
.PARAM R2 = 100
.PARAM G2 = {1/R2}
.PARAM GOUT = {1/ROUT}
.PARAM C2 = {1/(2*PI*R2*FPOLE2)}
.PARAM VDF = {VT*LOG(1 + IMAX/IS)}
IBIASM      INM 0  {IBIAS - IOFFS}
RINM      INM  8  {2*RINC}
RINP      INP  8  {2*RINC}
IBIAS       10 0   {IBIAS}
VOFFS       10 INP  {VOFFS}
EVP VPI 0 VP 0 1
EVM VMI 0 VM 0 1
VC          VPI 11  {VDROPOH + VDF}
VE          12 VMI  {VDROPOL + VDF}
D1          VM VP  D_1
RP          VP VM  15E3
ROUT        OUT 8  {ROUT}
GMO         8 OUT 9 8 {GOUT}
C2          9 8  {C2}
R2          9 8  {R2}
GM2         8 9 7 8 {G2}
RIN         INM 10  {RIN}
EGND        8  0  POLY(2) (VP,0) (VM,0) 0 .5 .5
D3         12 7  D_1
D2          7 11  D_1
C1          7 8  {C1}
R1          7 8  {R1}
GM1         8 7 VALUE = { LIMIT( GM1*V(10,INM), -IMAX, IMAX) }
.MODEL D_1 D( IS={IS} )
.ENDS

.SUBCKT idopamp In+ In- Out
+ Params: GAIN=1E12
EO         OUT 0  In+ In-  {GAIN}
.ENDS

.TEMP 27
.TRAN 4U 8M UIC
.OPTIONS ABSTOL=1U ITL2=20 TRTOL=7
.PROBE V(6)

V6          4 0 6.9
V5          0 11 6.9
V4          0 16 6.9
V3          17 0 6.9
V2          0 18 6.9
V1          19 0 6.9
Vin         10 0 DC 0 AC 1 0
+ PULSE ( 0 1 0 0 0 2M 4M )
R18         2 3 10K ; *DIST: UNIFORM 0 *
R17         3 1 10K ; *DIST: UNIFORM 0 *
XIOP1        0 3 1 IdOpamp
R16         4 5 1.51K ; *DIST: UNIFORM 0 *
R15         5 2 1K ; *DIST: UNIFORM 0 *
R14         6 5 1K ; *DIST: UNIFORM 0 *
XLM301A      0 5 2 IdOpamp
RES4        7 8 27K ; *DIST: NORMAL 0.1 *
R11         8 9 3K ; *DIST: UNIFORM 0 *
C2          7 8 100N ; *DIST: NORMAL 0.1 *
R12         10 7 10K ; *DIST: UNIFORM 0 *
XLM301A_2    0 7 8 IdOpamp
R10         11 9 3.7K ; *DIST: UNIFORM 0 *
R9          9 12 1K ; *DIST: UNIFORM 0 *
XLM301A_3    0 9 12 IdOpamp
QT1         14 6 13  Q_2N2222_N_1 
RES1        15 14 1K ; *DIST: UNIFORM 0 *
RES2        15 13 10K ; *DIST: NORMAL 0.1 *
C1          15 13 100N ; *DIST: NORMAL 0.1 *
XOP2         0 15 17 16 13 StdOpamp
+ PARAMS: GAIN=160K RIN=2MEG ROUT=75 SLEWRATE=10MEG FPOLE1=5 FPOLE2=1MEG VOFFS=2M IBIAS=70N IOFFS=3N VDROPOH=1.9 VDROPOL=1.9
XOP1         20 21 19 18 6 StdOpamp
+ PARAMS: GAIN=160K RIN=2MEG ROUT=75 SLEWRATE=10MEG FPOLE1=5 FPOLE2=1MEG VOFFS=2M IBIAS=70N IOFFS=3N VDROPOH=1.9 VDROPOL=1.9
R7          13 22 10K ; *DIST: UNIFORM 0 *
R8          22 23 10K ; *DIST: UNIFORM 0 *
XLM301A_4    0 22 23 IdOpamp
R6          10 15 1K ; *DIST: UNIFORM 0 *
R3          12 21 820 ; *DIST: UNIFORM 0 *
RES3        20 6 2.7K ; *DIST: UNIFORM 0 *
R1          23 20 1K ; *DIST: UNIFORM 0 *

.MODEL Q_2N2222_N_1 NPN( IS=11.9F NF=1 NR=1 RE=649M RC=1 
+      RB=10 VAF=56.7 VAR=28.3 ISE=146F ISC=146F 
+      ISS=0 NE=1.49 NC=1.49 NS=1 BF=215 
+      BR=5 IKF=143M IKR=143M CJC=13.1P CJE=30P 
+      CJS=0 VJC=2.87 VJE=500 VJS=750M MJC=330M 
+      MJE=100M MJS=0 TF=637P TR=82.8N EG=1.11 
+      KF=0 AF=1 )

.END