sum2 (PSpice format)
.SUBCKT IdOpamp In+ In- Out
+ Params: GAIN=1E12
*
EO         OUT 0  In+ In-  {GAIN}
.ENDS

.TEMP 27
.TRAN 2U 1M UIC
.DC LIN VG3 0 1 10M

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V(6,0)

VG3         1 7 DC 0 AC 1 0
+ PWL TIME_SCALE_FACTOR=250U VALUE_SCALE_FACTOR=500M
+      REPEAT FOREVER
+       (0, 0) (4U 1) (499.996M 1) (500.004M -1) (999.996M -1) (1,0) ENDREPEAT
VG3_DC      7 0 500M
VG2         2 8 DC 0 AC 1 0
+ PWL TIME_SCALE_FACTOR=500U VALUE_SCALE_FACTOR=500M
+      REPEAT FOREVER
+       (0, 0) (2U 1) (499.998M 1) (500.002M -1) (999.998M -1) (1,0) ENDREPEAT
VG2_DC      8 0 500M
VG1         3 9 DC 0 AC 1 0
+ PWL TIME_SCALE_FACTOR=1M VALUE_SCALE_FACTOR=500M
+      REPEAT FOREVER
+       (0, 0) (1U 1) (499.999M 1) (500.001M -1) (999.999M -1) (1,0) ENDREPEAT
VG1_DC      9 0 500M
XIOP1        4 5 6 IdOpamp
R5          5 0 1K 
R4          5 6 1K 
R3          3 4 1K 
R2          2 4 1K 
R1          1 4 1K 


.END
