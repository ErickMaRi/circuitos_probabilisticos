LINEAL (PSpice format)
.TEMP 27
.TRAN 20N 10U

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V(4,0)

VIN         3 0 DC 0 AC 1 0
+ PULSE ( 0 1 0  0  0  1e19 1e20 )
R2 1 0 1.0248774752379386K
L2 2 1 997.5829463226509u IC=0
R1 3 2 1.0126609095614814K
lin         4 3 1M IC=0 
C1 4 2 1.0186047034224694u

.END
