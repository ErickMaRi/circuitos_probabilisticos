PEAK DETECTOR
.TEMP 27
.TRAN 40N 20U

.OPTIONS ABSTOL=1U ITL1=150 ITL2=20 ITL4=2000 TRTOL=7 
.PROBE V([Vout])

V1          0 V- 2.5
Vin         5 0 DC 0 AC 1 0
+ SIN( 0 10M 500K 0 0 0 )
V1_2        V+ 0 2.5
XU2         3 Vout V+ V- Vout OPA354_0
XU1         5 6 V+ V- 7 OPA354_0
DSD1        7 3  D_BAT17_1 
R2          6 Vout 2K 
R1          8 3 3 
C2          6 7 5P IC=0 
C1          0 8 10N IC=0 

.MODEL D_BAT17_1 D( IS=139.7P N=1 BV=4 IBV=333N RS=13.22 
+      CJO=1P VJ=750M M=330M FC=500M TT=1.67N 
+      EG=1.11 XTI=3 KF=0 AF=1 )

* OPA354 SPICE MACRO-MODEL
*
*   REV. A    12 JANUARY 2004, BY W.K. SANDS
*
*   REV. B    4 JANUARY 2004 BY NEIL ALBAUGH: ADDED HEADER TEXT & EDITED TEXT
*
* THIS MACROMODEL HAS BEEN OPTIMIZED TO MODEL THE AC, DC, AND TRANSIENT RESPONSE PERFORMANCE WITHIN
*     THE DEVICE DATA SHEET SPECIFIED LIMITS.
*     CORRECT OPERATION OF THIS MACROMODEL HAS BEEN VERIFIED ON MICROSIM P-SPICE VER. 8.0 AND ON
*     PENZAR DEVELOPMENT TOPSPICE VER. 6.82D. FOR HELP WITH OTHER ANALOG SIMULATION SOFTWARE,
*     PLEASE CONSULT YOUR SOFTWARE SUPPLIER.
*
*
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
*
* BEGIN MODEL OPA354
*
* BEGIN NOTES
*
*
* MODEL TEMPERATURE RANGE IS -40 C TO +125 C, NOT ALL PARAMETERS ACCURATELY TRACK THOSE OF AN ACTUAL OPA357
* OVER THE FULL TEMPERATURE RANGE BUT ARE AS CLOSE AS PRACTICAL
*
* END NOTES
*
*
* BEGIN MODEL OPA354
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   4   5  2  1
.SUBCKT OPA354_0  3 4 5 2 1
* BEGIN SIMULATION NOTES
* FOR BEST RESULTS WHEN LOOKING AT INPUT BIAS CURRENTS
* SET ABSTOL FROM 1E-13 TO 3E-13
* FOR AID IN DC CONVERGENCE SET ITL1 FROM 400 TO 4000
* FOR AID IN TRANSIENT ANALYSIS SET ITL4 FROM 50 TO 500
* MODEL TEMPERATURE RANGE IS
* -40 C TO +125 C, NOT ALL
* PARAMETERS TRACK THOSE OF
* THE REAL PART VS TEMPERATURE
* END SIMULATION NOTES
* BEGIN MODEL FEATURES
* OPEN LOOP GAIN AND PHASE
* INPUT OFFSET VOLTAGE CHANGE AT THE
* RAIL-TO-RAIL INPUT TRANSITION POINT
* INPUT VOLTAGE NOISE WITH 1/F
* INPUT CURRENT NOISE
* INPUT BIAS CURRENT
* INPUT CAPACITANCE
* INPUT COMMON MODE VOLTAGE RANGE
* INPUT CLAMPS TO RAILS
* CMRR WITH FREQUENCY EFFECTS
* PSRR WITH FREQUENCY EFFECTS
* SLEW RATE
* QUIESCENT CURRENT
* RAIL TO RAIL OUTPUT STAGE
* HIGH CLOAD EFFECTS
* CLASS AB BIAS IN OUTPUT STAGE
* OUTPUT CURRENT THROUGH SUPPLIES
* OUTPUT CURRENT LIMITING
* OUTPUT CLAMPS TO RAILS
* OUTPUT SWING VS OUTPUT CURRENT
* END MODEL FEATURES
Q20 6 7 8 QLN
R3 9 10 20
R4 11 10 20
R10 7 12 1E3
R11 13 14 1E3
R12 14 5 2.5
R13 2 12 2.5
R16 15 16 1E3
R17 17 18 2.5
R18 8 19 2.5
D5 20 5 DD
D6 2 20 DD
D7 21 0 DIN
D8 22 0 DIN
I8 0 21 0.1E-3
I9 0 22 0.1E-3
E2 8 0 2 0 1
E3 18 0 5 0 1
D9 23 0 DVN
D10 24 0 DVN
I10 0 23 0.1E-3
I11 0 24 0.1E-3
E4 25 4 23 24 0.18
G2 26 4 21 22 5E-7
R22 2 5 100E6
E5 27 0 18 0 1
E6 28 0 8 0 1
E7 29 0 30 0 1
R30 27 31 1E4
R31 28 32 1E5
R32 29 33 1E5
R33 0 31 1
R34 0 32 10
R35 0 33 10
E10 34 3 33 0 0.4
R36 35 30 1K
R37 30 36 1K
C6 27 31 0.2E-12
C7 28 32 100E-12
C8 29 33 2E-12
E11 37 34 32 0 0.5
E12 26 37 31 0 3.3
E14 38 8 18 8 0.5
D11 15 18 DD
D12 8 15 DD
M1 39 40 12 12 NOUT L=3U W=800U
M2 41 42 14 14 POUT L=3U W=800U
M3 43 43 17 17 POUT L=3U W=800U
M4 44 45 9 9 PIN L=3U W=160U
M5 46 25 11 11 PIN L=3U W=160U
M8 47 47 19 19 NOUT L=3U W=800U
R43 48 42 100
R44 49 40 100
G3 15 38 50 38 0.2E-3
R45 38 15 200E6
C12 16 20 1E-12
R46 8 44 2E3
R47 8 46 2E3
C13 44 46 0.125E-12
C14 26 0 0.68E-12
C15 25 0 0.68E-12
C16 20 0 0.5E-12
D13 40 6 DD
D14 51 42 DD
Q15 51 13 18 QLP
V18 26 45 0.7E-3
M16 52 53 54 54 NIN L=3U W=160U
R53 55 54 20
M17 56 25 57 57 NIN L=3U W=160U
R54 55 57 20
R55 52 18 2E3
R56 56 18 2E3
C20 52 56 0.125E-12
V19 45 53 -2E-3
M18 58 59 60 60 PIN L=6U W=500U
M19 61 62 18 18 PIN L=6U W=500U
V20 18 59 1.3
M21 55 58 8 8 NIN L=6U W=500U
M22 58 58 8 8 NIN L=6U W=500U
G6 15 38 63 38 0.2E-3
E17 36 0 26 0 1
E18 35 0 4 0 1
M23 62 62 18 18 PIN L=6U W=500U
V21 61 10 0
R59 20 41 5
R60 39 20 5
J1 64 26 64 JNC
J2 64 25 64 JNC
J3 25 65 25 JNC
J4 26 65 26 JNC
C21 26 25 0.5E-12
E19 66 38 56 52 1
R61 66 63 1E4
C22 63 38 0.125E-12
E20 67 38 46 44 1
R62 67 50 1E4
C23 50 38 0.125E-12
G7 68 38 15 38 -1E-3
G8 38 69 15 38 1E-3
G9 38 70 47 8 1E-3
G10 71 38 18 43 1E-3
D17 71 68 DD
D18 69 70 DD
R66 68 71 100E6
R67 70 69 100E6
R68 71 18 1E3
R69 8 70 1E3
E23 18 48 18 71 1
E24 49 8 70 8 1
R70 69 38 1E6
R71 70 38 1E6
R72 38 71 1E6
R73 38 68 1E6
G11 5 2 72 0 3.55E-3
R75 37 26 1E9
R76 34 37 1E9
R77 3 34 1E9
R78 4 25 1E9
R79 38 50 1E9
R80 38 63 1E9
R81 48 18 1E9
R82 8 49 1E9
R83 30 0 1E9
R85 60 61 1E3
G14 62 8 73 0 400E-6
G15 43 47 73 0 1.35E-3
E48 74 15 73 0 30
E49 75 38 73 0 -30
V49 76 75 15
V50 77 74 -15
R127 74 0 1E12
R128 75 0 1E12
M41 38 77 15 78 PSW L=1.5U W=150U
M42 15 76 38 79 NSW L=1.5U
R129 78 0 1E12
R130 79 0 1E12
M43 80 81 8 8 NEN L=3U W=300U
M44 82 80 8 8 NEN L=3U W=3000U
R131 80 18 1E4
R132 82 83 1E6
V51 83 8 1
M45 84 84 18 18 PEN L=6U W=60U
M46 81 84 18 18 PEN L=6U W=60U
I20 84 8 0.2E-6
C26 81 0 1E-12
E50 73 0 85 8 1
V52 82 85 1.111E-6
R133 8 85 1E12
C32 18 80 15E-12
C33 83 82 0.15E-12
I21 5 2 3.4E-6
L1 20 1 4E-9
R150 20 1 400
V78 18 64 0
V79 65 8 0
I22 25 0 1E-12
I23 26 0 1E-12
M47 86 80 8 8 NEN L=3U W=3000U
R152 86 83 1E6
C34 83 86 0.005E-12
V80 86 87 1.111E-6
R153 8 87 1E12
E53 72 0 87 8 1
R154 0 72 1E12
R155 43 18 1E9
R156 8 47 1E9
R157 12 40 1E9
R158 14 42 1E9
R159 81 18 10E6
RG1 73 0 1E9
.MODEL DVN D KF=8E-12 IS=1E-16
.MODEL DD D
.MODEL DIN D
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL JNC NJF
.MODEL POUT PMOS KP=200U VTO=-0.7
.MODEL NOUT NMOS KP=200U VTO=0.7
.MODEL PIN PMOS KP=200U VTO=-0.7
.MODEL NIN NMOS KP=200U VTO=0.7
.MODEL NEN NMOS KP=200U VTO=0.5 IS=1E-18
.MODEL PEN PMOS KP=200U VTO=-0.7 IS=1E-18
.MODEL PSW PMOS KP=200U VTO=-7.5 IS=1E-18
.MODEL NSW NMOS KP=200U VTO=7.5 IS=1E-18
.ENDS


.END
