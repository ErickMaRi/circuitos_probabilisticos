sum (PSpice format)
.SUBCKT STDOPAMP  INP INM VP VM OUT
+ PARAMS: GAIN=200K RIN=2MEG RINC=1E9 ROUT=75 SLEWRATE=500K FPOLE1=5 FPOLE2=1MEG 
+         VDROPOH=1.9 VDROPOL=1.9 VOFFS=1M IBIAS=80N IOFFS=20N 
.PARAM PI = 3.141592
.PARAM IS = 1.0E-12
.PARAM VT = 0.02585
.PARAM IMAX = 100.0E-2
.PARAM C1 = {IMAX/SLEWRATE}
.PARAM R1 = {1/(2*PI*C1*FPOLE1)}
.PARAM GM1 = {GAIN/R1}
.PARAM R2 = 100
.PARAM G2 = {1/R2}
.PARAM GOUT = {1/ROUT}
.PARAM C2 = {1/(2*PI*R2*FPOLE2)}
.PARAM VDF = {VT*LOG(1 + IMAX/IS)}
IBIASM      INM 0  {IBIAS - IOFFS}
RINM      INM  8  {2*RINC}
RINP      INP  8  {2*RINC}
IBIAS       10 0   {IBIAS}
VOFFS       10 INP  {VOFFS}
EVP VPI 0 VP 0 1
EVM VMI 0 VM 0 1
VC          VPI 11  {VDROPOH + VDF}
VE          12 VMI  {VDROPOL + VDF}
D1          VM VP  D_1
RP          VP VM  15E3
ROUT        OUT 8  {ROUT}
GMO         8 OUT 9 8 {GOUT}
C2          9 8  {C2}
R2          9 8  {R2}
GM2         8 9 7 8 {G2}
RIN         INM 10  {RIN}
EGND        8  0  POLY(2) (VP,0) (VM,0) 0 .5 .5
D3         12 7  D_1
D2          7 11  D_1
C1          7 8  {C1}
R1          7 8  {R1}
GM1         8 7 VALUE = { LIMIT( GM1*V(10,INM), -IMAX, IMAX) }
.MODEL D_1 D( IS={IS} )
.ENDS

.TEMP 27
.AC DEC 20 10 1MEG
.TRAN 2N 1U 0

.OPTIONS ABSTOL=1P ITL1=150 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V(4,0)

VS5         1 0 5
VS4         2 0 5
VS3         3 0 5
VS2         0 5 5
VS1         6 0 5
R5          7 0 1K 
R4          7 4 1K 
R3          3 8 1K 
R2          2 8 1K 
R1          1 8 1K 
XOP1         8 7 6 5 4 StdOpamp
+ PARAMS: GAIN=160K RIN=2MEG ROUT=50 SLEWRATE=70MEG FPOLE1=75 FPOLE2=4.7MEG VOFFS=4M IBIAS=150N IOFFS=30N VDROPOH=2 VDROPOL=2


.END
