10MHZ_ACTIVE_LPF_FOR_PSPICE (PSpice format)
.TEMP 27
.TRAN 4N 2U

.OPTIONS ABSTOL=1U ITL1=100 ITL2=20 ITL4=10 TRTOL=7 
.PROBE V(140, 0)

Vbias       0 4 -2.5
Vin         5 131 DC 0 AC 1 0
+ SIN( 0 1 1MEG 0 0 0 )
Vin_DC      131 4 -2.5
V1          2 0 5
XU1         0 1 2 0 140 OPA380_0
C2          6 0 47P IC=0 
R3          5 6 576 
R2          6 1 1.37K 
R1          6 140 576 
C1          1 140 6.8P IC=0 


* OPA380 SPICE MACRO-MODEL 
*          
*   REV. A    26 MARCH 2004, BY W.K. SANDS
*
*   REV. B    2 APRIL 2004 BY NEIL ALBAUGH: ADDED HEADER TEXT & EDITED TEXT
*
* THIS MACROMODEL HAS BEEN OPTIMIZED TO MODEL THE AC, DC, AND TRANSIENT RESPONSE PERFORMANCE WITHIN 
*     THE DEVICE DATA SHEET SPECIFIED LIMITS. 
*     CORRECT OPERATION OF THIS MACROMODEL HAS BEEN VERIFIED ON MICROSIM P-SPICE VER. 8.0 AND ON 
*     PENZAR DEVELOPMENT TOPSPICE VER. 6.82D. FOR HELP WITH OTHER ANALOG SIMULATION SOFTWARE, 
*     PLEASE CONSULT YOUR SOFTWARE SUPPLIER. 
*
*  
* ------------------------------------------------------------------------
*|(C) COPYRIGHT TEXAS INSTRUMENTS INCORPORATED 2007. ALL RIGHTS RESERVED. |
*|                                                                        |
*|THIS MODEL IS DESIGNED AS AN AID FOR CUSTOMERS OF TEXAS INSTRUMENTS.    |
*|NO WARRANTIES, EITHER EXPRESSED OR IMPLIED, WITH RESPECT TO THIS MODEL  |
*|OR ITS FITNESS FOR A PARTICULAR PURPOSE IS CLAIMED BY TEXAS INSTRUMENTS |
*|OR THE AUTHOR.  THE MODEL IS LICENSED SOLELY ON AN "AS IS" BASIS.  THE  |
*|ENTIRE RISK AS TO ITS QUALITY AND PERFORMANCE IS WITH THE CUSTOMER.     |
* ------------------------------------------------------------------------
*
*
* BEGIN NOTES
*
*
* MODEL TEMPERATURE RANGE IS -40 C TO +125 C, NOT ALL PARAMETERS ACCURATELY TRACK THOSE OF AN ACTUAL OPA380 
* OVER THE FULL TEMPERATURE RANGE BUT ARE AS CLOSE AS PRACTICAL
*
* CMRR ACCURACY AT DC HAS BEEN TRADED OFF FOR IMPROVED CONVERGENCE - 
* MODELED CMRR DC IS ONLY 86 DB; ACTUAL OPA380 IS MUCH HIGHER
*
* END NOTES
*
* BEGIN FEATURES
*
* OPEN LOOP GAIN AND PHASE
* INPUT OFFSET VOLTAGE
* TEMPERATURE EFFECTS SAME
* INPUT VOLTAGE NOISE
* INPUT CURRENT NOISE
* INPUT BIAS CURRENT
* TEMPERATURE EFFECTS SAME
* INPUT CAPACITANCE
* INPUT COMMON MODE VOLTAGE RANGE
* INPUT CLAMPS TO RAILS
* CMRR WITH FREQUENCY EFFECTS
* PSRR WITH FREQUENCY EFFECTS
* SLEW RATE
* QUIESCENT CURRENT
* QUIESCENT CURRENT VS VOLTAGE
* RAIL TO RAIL OUTPUT STAGE
* HIGH CLOAD EFFECTS
* CLASS AB BIAS IN OUTPUT STAGE
* OUTPUT CURRENT THROUGH SUPPLIES
* OUTPUT CURRENT LIMITING
* OUTPUT CLAMPS TO RAILS
* OUTPUT SWING VS OUTPUT CURRENT
* OUTPUT WILL SWING SLIGHTLY
* BELOW -V W EXTERNAL PULLDOWN
* TO A SUPPLY MORE NEGATIVE
* THAN -V
* END FEATURES
*
* BEGIN MODEL OPA380
*
* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER  3   2   1  4  6
.SUBCKT OPA380_0  3 2 1 4 6
*
R81 10 1 1
R82 4 11 1
R84 12 13 700
R85 14 15 1
R86 16 17 1
D21 9 1 DD
D22 4 9 DD
D23 18 0 DIN
D24 19 0 DIN
I24 0 18 0.1E-3
I25 0 19 0.1E-3
E25 16 0 4 0 1
E26 15 0 1 0 1
G13 20 21 18 19 5E-6
E28 22 0 15 0 1
E29 23 0 16 0 1
E30 24 0 25 0 1
R88 22 26 1E6
R89 23 27 1E6
R90 24 28 1E6
R91 0 26 100
R92 0 27 100
R93 0 28 100
E31 29 3 28 0 9.5E-4
R94 30 25 1E3
R95 25 31 1E3
C29 22 26 0.2E-12
C30 23 27 0.2E-12
C31 24 28 6E-9
E32 32 29 27 0 0.042
E33 33 32 26 0 0.002
E34 34 16 15 16 0.5
D27 12 15 DD
D28 16 12 DD
M24 35 36 11 11 NOUT L=3U W=4000U
M25 37 38 10 10 POUT L=3U W=4000U
M26 39 39 14 14 POUT L=3U W=4000U
M27 40 41 42 42 PIN L=3U W=40U
M28 43 44 42 42 PIN L=3U W=40U
M29 45 45 17 17 NOUT L=3U W=4000U
R96 46 38 100
R97 47 36 100
G14 12 34 48 34 0.2E-3
R98 34 12 100E3
C32 13 9 27E-12
R99 16 40 6E3
R100 16 43 6E3
C33 40 43 3E-12
C34 20 0 1E-12
C35 21 0 1E-12
C36 9 0 1E-12
V27 20 49 -10E-6
M33 50 51 15 15 PIN L=6U W=500U
E35 31 0 20 0 1
E36 30 0 21 0 1
M36 51 51 15 15 PIN L=6U W=500U
V30 50 42 0.8
R105 9 37 40
R106 35 9 22
J5 52 20 52 JC
J6 52 21 52 JC
J7 21 53 21 JC
J8 20 53 20 JC
E38 54 34 43 40 1
R108 54 48 10E3
C40 48 34 1.5E-12
G16 55 34 12 34 -1E-3
G17 34 56 12 34 1E-3
G18 34 57 45 16 1E-3
G19 58 34 15 39 1E-3
D31 58 55 DD
D32 56 57 DD
R110 55 58 100E6
R111 57 56 100E6
R112 58 15 1E3
R113 16 57 1E3
E39 15 46 15 58 1
E40 47 16 57 16 1
R114 56 34 1E6
R115 57 34 1E6
R116 34 58 1E6
R117 34 55 1E6
C46 59 20 0.1E-12
R122 0 59 220
E41 59 0 18 19 210
V45 15 52 0.2
V46 53 16 0.2
E56 20 33 60 0 30E-6
D51 61 0 DD
R139 0 60 1E9
R140 0 61 1E9
V55 61 60 0.65
I35 0 61 1E-3
R141 49 41 84E3
R142 44 21 84E3
C49 20 21 1E-12
Q23 62 63 64 QLN
R150 63 65 1E3
R151 66 67 1E3
R152 68 1 2
R153 4 69 2
R155 70 71 680
R156 72 73 2
R157 64 74 2
D54 75 1 DD
D55 4 75 DD
D56 76 0 DIN
D57 77 0 DIN
I36 0 76 0.1E-3
I37 0 77 0.1E-3
E57 64 0 4 0 1
E58 73 0 1 0 1
D58 78 0 DVN
D59 79 0 DVN
I38 0 78 0.1E-3
I39 0 79 0.1E-3
E59 80 2 78 79 0.025
G24 81 2 76 77 1.6E-6
R158 4 1 2E3
E60 82 0 73 0 1
E61 83 0 64 0 1
E62 84 0 85 0 1
R160 82 86 1E4
R161 83 87 1E5
R162 84 88 1E5
R163 0 86 1
R164 0 87 10
R165 0 88 10
E63 89 90 88 0 0.03
R166 91 85 1E3
R167 85 92 1E3
C51 82 86 10E-12
C52 83 87 10E-12
C53 84 88 10E-12
E64 93 89 87 0 0.3
E65 81 93 86 0 0.3
E66 94 64 73 64 0.5
D60 70 73 DD
D61 64 70 DD
M52 95 96 69 69 NOUT L=3U W=450U
M53 97 98 68 68 POUT L=3U W=950U
M54 99 99 72 72 POUT L=3U W=950U
M55 100 101 102 102 PIN L=3U W=270U
M56 103 104 102 102 PIN L=3U W=270U
M57 105 105 74 74 NOUT L=3U W=450U
R168 106 98 100
R169 107 96 100
G25 70 94 108 94 0.2E-3
R170 94 70 2E6
C54 71 75 1.65E-12
R171 64 100 2E3
R172 64 103 2E3
C55 100 103 0.11E-12
C56 81 0 3E-12
C57 80 0 3E-12
C58 75 0 0.5E-12
D62 96 62 DD
D63 109 98 DD
Q24 109 67 73 QLP
V58 81 110 0
M58 111 112 73 73 PIN L=6U W=500U
E67 92 0 81 0 1
E68 91 0 2 0 1
M59 112 112 73 73 PIN L=6U W=500U
V59 111 102 1
R173 113 97 0.25
R174 95 75 4
J11 114 81 114 JNC
J12 114 80 114 JNC
J13 80 115 80 JNC
J14 81 115 81 JNC
C59 81 116 1.1E-12
E69 117 94 103 100 1
R175 117 108 1E4
C60 108 94 0.11E-12
G26 118 94 70 94 -1E-3
G27 94 119 70 94 1E-3
G28 94 120 105 64 1E-3
G29 121 94 73 99 1E-3
D64 121 118 DD
D65 119 120 DD
R176 118 121 100E6
R177 120 119 100E6
R178 121 73 1E3
R179 64 120 1E3
E70 73 106 73 121 1
E71 107 64 120 64 1
R180 119 94 1E6
R181 120 94 1E6
R182 94 121 1E6
R183 94 118 1E6
R184 93 81 1E9
R185 89 93 1E9
R186 90 89 1E9
R187 2 80 1E9
R188 94 108 1E9
R189 106 73 1E9
R190 64 107 1E9
R191 85 0 1E9
I41 1 4 1.5E-3
L2 75 6 4E-9
R200 75 6 400
V79 73 114 0
V80 115 64 0
R204 99 73 1E8
R205 64 105 1E8
R206 69 96 1E8
R207 68 98 1E8
R209 116 80 100
R226 104 80 400
R227 101 110 400
E96 73 66 1 68 1
E97 65 64 69 4 1
R314 112 73 1E9
R316 9 122 100E3
C69 122 3 75E-12
C70 21 9 67E-12
R318 123 21 900E3
R320 2 123 100E3
C72 123 6 115E-15
V118 113 75 0.4
R325 20 33 1E9
R326 32 33 1E9
R327 29 32 1E9
R328 3 29 1E9
I49 99 105 2E-3
I50 112 64 360E-6
I51 51 16 37.5E-6
I52 39 45 20E-6
C74 59 21 0.1E-12
G36 80 0 124 0 10E-12
I53 80 0 3E-12
I54 0 125 1E-3
D67 125 0 DD
V120 125 126 0.7
R329 0 126 1E6
E98 127 0 126 0 -571
R330 0 127 1E6
R331 128 127 1E3
G37 20 0 124 0 10E-12
I55 20 0 3E-12
R332 0 129 1E6
V121 130 0 73.5
D68 131 129 DD
D69 128 129 DD
R333 131 130 1E3
V122 129 132 72.8
R334 0 132 1E6
E99 124 0 132 0 1.5
R335 0 124 1E6
V123 90 122 -15E-3
R338 39 15 1E9
R339 16 45 1E9
R340 11 36 1E9
R341 10 38 1E9
R343 51 15 1E9
R344 34 9 100E3
R345 94 75 50E3
.MODEL DVN D KF=2E-11 IS=1E-16
.MODEL DD D
.MODEL DIN D
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL JNC NJF
.MODEL JC NJF IS=1E-18
.MODEL JE NJF IS=1E-17
.MODEL POUT PMOS KP=200U VTO=-0.7
.MODEL NOUT NMOS KP=200U VTO=0.7
.MODEL PIN PMOS KP=200U VTO=-0.7
.MODEL NIN NMOS KP=200U VTO=0.7
.ENDS


.END
